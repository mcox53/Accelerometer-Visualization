-- Author: M. Cox
-- Date: 11/6/18
-- Description: Converts the desired PWM frequency to an evenly spaced 8 bit address.
-- The generated address will be used for the given Sine wave LUT

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity freq_to_addr_LUT is 
	port(
		freq 	: in std_logic_vector(13 downto 0);
		addr	: out std_logic_vector(7 downto 0)
		);
end freq_to_addr_LUT;

architecture behavioral of freq_to_addr_LUT is

begin
	with freq select
		addr <= X"00" when "00000000000000",
				X"00" when "00000001000000",
				X"01" when "00000010000000",
				X"02" when "00000011000000",
				X"02" when "00000100000000",
				X"03" when "00000101000000",
				X"04" when "00000110000000",
				X"04" when "00000111000000",
				X"05" when "00001000000000",
				X"06" when "00001001000000",
				X"06" when "00001010000000",
				X"07" when "00001011000000",
				X"08" when "00001100000000",
				X"08" when "00001101000000",
				X"09" when "00001110000000",
				X"0a" when "00001111000000",
				X"0a" when "00010000000000",
				X"0b" when "00010001000000",
				X"0c" when "00010010000000",
				X"0c" when "00010011000000",
				X"0d" when "00010100000000",
				X"0e" when "00010101000000",
				X"0e" when "00010110000000",
				X"0f" when "00010111000000",
				X"10" when "00011000000000",
				X"10" when "00011001000000",
				X"11" when "00011010000000",
				X"12" when "00011011000000",
				X"12" when "00011100000000",
				X"13" when "00011101000000",
				X"14" when "00011110000000",
				X"14" when "00011111000000",
				X"15" when "00100000000000",
				X"16" when "00100001000000",
				X"16" when "00100010000000",
				X"17" when "00100011000000",
				X"18" when "00100100000000",
				X"18" when "00100101000000",
				X"19" when "00100110000000",
				X"1a" when "00100111000000",
				X"1a" when "00101000000000",
				X"1b" when "00101001000000",
				X"1c" when "00101010000000",
				X"1c" when "00101011000000",
				X"1d" when "00101100000000",
				X"1e" when "00101101000000",
				X"1e" when "00101110000000",
				X"1f" when "00101111000000",
				X"20" when "00110000000000",
				X"21" when "00110001000000",
				X"21" when "00110010000000",
				X"22" when "00110011000000",
				X"23" when "00110100000000",
				X"23" when "00110101000000",
				X"24" when "00110110000000",
				X"25" when "00110111000000",
				X"25" when "00111000000000",
				X"26" when "00111001000000",
				X"27" when "00111010000000",
				X"27" when "00111011000000",
				X"28" when "00111100000000",
				X"29" when "00111101000000",
				X"29" when "00111110000000",
				X"2a" when "00111111000000",
				X"2b" when "01000000000000",
				X"2b" when "01000001000000",
				X"2c" when "01000010000000",
				X"2d" when "01000011000000",
				X"2d" when "01000100000000",
				X"2e" when "01000101000000",
				X"2f" when "01000110000000",
				X"2f" when "01000111000000",
				X"30" when "01001000000000",
				X"31" when "01001001000000",
				X"31" when "01001010000000",
				X"32" when "01001011000000",
				X"33" when "01001100000000",
				X"33" when "01001101000000",
				X"34" when "01001110000000",
				X"35" when "01001111000000",
				X"35" when "01010000000000",
				X"36" when "01010001000000",
				X"37" when "01010010000000",
				X"37" when "01010011000000",
				X"38" when "01010100000000",
				X"39" when "01010101000000",
				X"39" when "01010110000000",
				X"3a" when "01010111000000",
				X"3b" when "01011000000000",
				X"3b" when "01011001000000",
				X"3c" when "01011010000000",
				X"3d" when "01011011000000",
				X"3d" when "01011100000000",
				X"3e" when "01011101000000",
				X"3f" when "01011110000000",
				X"40" when "01011111000000",
				X"40" when "01100000000000",
				X"41" when "01100001000000",
				X"42" when "01100010000000",
				X"42" when "01100011000000",
				X"43" when "01100100000000",
				X"44" when "01100101000000",
				X"44" when "01100110000000",
				X"45" when "01100111000000",
				X"46" when "01101000000000",
				X"46" when "01101001000000",
				X"47" when "01101010000000",
				X"48" when "01101011000000",
				X"48" when "01101100000000",
				X"49" when "01101101000000",
				X"4a" when "01101110000000",
				X"4a" when "01101111000000",
				X"4b" when "01110000000000",
				X"4c" when "01110001000000",
				X"4c" when "01110010000000",
				X"4d" when "01110011000000",
				X"4e" when "01110100000000",
				X"4e" when "01110101000000",
				X"4f" when "01110110000000",
				X"50" when "01110111000000",
				X"50" when "01111000000000",
				X"51" when "01111001000000",
				X"52" when "01111010000000",
				X"52" when "01111011000000",
				X"53" when "01111100000000",
				X"54" when "01111101000000",
				X"54" when "01111110000000",
				X"55" when "01111111000000",
				X"56" when "10000000000000",
				X"56" when "10000001000000",
				X"57" when "10000010000000",
				X"58" when "10000011000000",
				X"58" when "10000100000000",
				X"59" when "10000101000000",
				X"5a" when "10000110000000",
				X"5a" when "10000111000000",
				X"5b" when "10001000000000",
				X"5c" when "10001001000000",
				X"5c" when "10001010000000",
				X"5d" when "10001011000000",
				X"5e" when "10001100000000",
				X"5e" when "10001101000000",
				X"5f" when "10001110000000",
				X"60" when "10001111000000",
				X"61" when "10010000000000",
				X"61" when "10010001000000",
				X"62" when "10010010000000",
				X"63" when "10010011000000",
				X"63" when "10010100000000",
				X"64" when "10010101000000",
				X"65" when "10010110000000",
				X"65" when "10010111000000",
				X"66" when "10011000000000",
				X"67" when "10011001000000",
				X"67" when "10011010000000",
				X"68" when "10011011000000",
				X"69" when "10011100000000",
				X"69" when "10011101000000",
				X"6a" when "10011110000000",
				X"6b" when "10011111000000",
				X"6b" when "10100000000000",
				X"6c" when "10100001000000",
				X"6d" when "10100010000000",
				X"6d" when "10100011000000",
				X"6e" when "10100100000000",
				X"6f" when "10100101000000",
				X"6f" when "10100110000000",
				X"70" when "10100111000000",
				X"71" when "10101000000000",
				X"71" when "10101001000000",
				X"72" when "10101010000000",
				X"73" when "10101011000000",
				X"73" when "10101100000000",
				X"74" when "10101101000000",
				X"75" when "10101110000000",
				X"75" when "10101111000000",
				X"76" when "10110000000000",
				X"77" when "10110001000000",
				X"77" when "10110010000000",
				X"78" when "10110011000000",
				X"79" when "10110100000000",
				X"79" when "10110101000000",
				X"7a" when "10110110000000",
				X"7b" when "10110111000000",
				X"7b" when "10111000000000",
				X"7c" when "10111001000000",
				X"7d" when "10111010000000",
				X"7d" when "10111011000000",
				X"7e" when "10111100000000",
				X"7f" when "10111101000000",
				X"80" when "10111110000000",
				X"80" when "10111111000000",
				X"81" when "11000000000000",
				X"82" when "11000001000000",
				X"82" when "11000010000000",
				X"83" when "11000011000000",
				X"84" when "11000100000000",
				X"84" when "11000101000000",
				X"85" when "11000110000000",
				X"86" when "11000111000000",
				X"86" when "11001000000000",
				X"87" when "11001001000000",
				X"88" when "11001010000000",
				X"88" when "11001011000000",
				X"89" when "11001100000000",
				X"8a" when "11001101000000",
				X"8a" when "11001110000000",
				X"8b" when "11001111000000",
				X"8c" when "11010000000000",
				X"8c" when "11010001000000",
				X"8d" when "11010010000000",
				X"8e" when "11010011000000",
				X"8e" when "11010100000000",
				X"8f" when "11010101000000",
				X"90" when "11010110000000",
				X"90" when "11010111000000",
				X"91" when "11011000000000",
				X"92" when "11011001000000",
				X"92" when "11011010000000",
				X"93" when "11011011000000",
				X"94" when "11011100000000",
				X"94" when "11011101000000",
				X"95" when "11011110000000",
				X"96" when "11011111000000",
				X"96" when "11100000000000",
				X"97" when "11100001000000",
				X"98" when "11100010000000",
				X"98" when "11100011000000",
				X"99" when "11100100000000",
				X"9a" when "11100101000000",
				X"9a" when "11100110000000",
				X"9b" when "11100111000000",
				X"9c" when "11101000000000",
				X"9c" when "11101001000000",
				X"9d" when "11101010000000",
				X"9e" when "11101011000000",
				X"9e" when "11101100000000",
				X"9f" when "11101101000000",
				X"a0" when "11101110000000",
				X"a1" when "11101111000000",
				X"a1" when "11110000000000",
				X"a2" when "11110001000000",
				X"a3" when "11110010000000",
				X"a3" when "11110011000000",
				X"a4" when "11110100000000",
				X"a5" when "11110101000000",
				X"a5" when "11110110000000",
				X"a6" when "11110111000000",
				X"a7" when "11111000000000",
				X"a7" when "11111001000000",
				X"a8" when "11111010000000",
				X"a9" when "11111011000000",
				X"a9" when "11111100000000",
				X"aa" when "11111101000000",
				X"ab" when "11111110000000",
				X"ab" when "11111111000000",
				X"00" when others;
end behavioral;